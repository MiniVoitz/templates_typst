module foo (
  input logic [13:0] a
);

endmodule